// megafunction wizard: %LPM_LATCH%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: lpm_latch 

// ============================================================
// File Name: ADD_LATCH.v
// Megafunction Name(s):
// 			lpm_latch
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 9.0 Build 132 02/25/2009 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2009 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module ADD_LATCH (
	aset,
	data,
	gate,
	q);

	input	  aset;
	input	[5:0]  data;
	input	  gate;
	output	[5:0]  q;

	wire [5:0] sub_wire0;
	wire [5:0] q = sub_wire0[5:0];

	lpm_latch	lpm_latch_component (
				.data (data),
				.gate (gate),
				.aset (aset),
				.q (sub_wire0),
				.aclr (1'b0),
				.aconst (1'b0));
	defparam
		lpm_latch_component.lpm_type = "LPM_LATCH",
		lpm_latch_component.lpm_width = 6;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: aclr NUMERIC "0"
// Retrieval info: PRIVATE: aset NUMERIC "1"
// Retrieval info: PRIVATE: nBit NUMERIC "6"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_LATCH"
// Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "6"
// Retrieval info: USED_PORT: aset 0 0 0 0 INPUT NODEFVAL aset
// Retrieval info: USED_PORT: data 0 0 6 0 INPUT NODEFVAL data[5..0]
// Retrieval info: USED_PORT: gate 0 0 0 0 INPUT NODEFVAL gate
// Retrieval info: USED_PORT: q 0 0 6 0 OUTPUT NODEFVAL q[5..0]
// Retrieval info: CONNECT: @data 0 0 6 0 data 0 0 6 0
// Retrieval info: CONNECT: q 0 0 6 0 @q 0 0 6 0
// Retrieval info: CONNECT: @gate 0 0 0 0 gate 0 0 0 0
// Retrieval info: CONNECT: @aset 0 0 0 0 aset 0 0 0 0
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: GEN_FILE: TYPE_NORMAL ADD_LATCH.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL ADD_LATCH.inc TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL ADD_LATCH.cmp TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL ADD_LATCH.bsf TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL ADD_LATCH_inst.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL ADD_LATCH_bb.v TRUE
// Retrieval info: LIB_FILE: lpm
