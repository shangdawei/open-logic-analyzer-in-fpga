module TestOutput(ain,bin,cin,out,Allout);

	input ain;
	input bin;
	input cin;
	output out;
	output [14:0] Allout;

	assign	out=(ain && bin) || cin;
	assign	Allout[0]=ain;
	assign	Allout[1]=ain;
	assign	Allout[2]=ain;
	assign	Allout[3]=ain;
	assign	Allout[4]=bin;
	assign	Allout[5]=bin;
	assign	Allout[6]=bin;
	assign	Allout[7]=bin;
	assign	Allout[8]=cin;
	assign	Allout[9]=cin;
	assign	Allout[10]=cin;
	assign	Allout[11]=cin;
	assign	Allout[12]=out;
	assign	Allout[13]=out;
	assign	Allout[14]=out;

endmodule
